library verilog;
use verilog.vl_types.all;
entity TB_EQU_SOLVER is
end TB_EQU_SOLVER;
